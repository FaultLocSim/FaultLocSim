module test;
reg a[];
reg b[];
initial begin
b = new[3];
end
endmodule
