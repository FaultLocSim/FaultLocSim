module a(
    a,
);
endmodule
