module test();

function void do_nothing();
  ;
endfunction

initial do_nothing();

endmodule
