module top;
    wire [3:0][2:0] arr;
    assign arr[2+:2] = 1;
endmodule
