module top;

a b (
    .*
);

endmodule
